// Verilog test fixture created from schematic C:\Xilinx\Lab1\Lab_3part2\zrodlo.sch - Fri Apr 17 21:05:17 2020

`timescale 1ns / 1ps

module zrodlo_zrodlo_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   zrodlo UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
