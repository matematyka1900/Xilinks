`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:24:28 04/24/2020 
// Design Name: 
// Module Name:    modul 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module modul(
	input [1:0] a,
	input [1:0] b,
	output [2:0] y
    );
	assign y = a + b;

endmodule
