// Verilog test fixture created from schematic C:\Xilinx\lab_3part4\schema.sch - Sat Apr 18 00:22:02 2020

`timescale 1ns / 1ps

module schema_schema_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   schema UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
